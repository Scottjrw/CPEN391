
module test_pixel_cluster_qsys (
	clk_clk,
	reset_reset_n,
	pixel_cluster_leds);	

	input		clk_clk;
	input		reset_reset_n;
	output	[9:0]	pixel_cluster_leds;
endmodule
