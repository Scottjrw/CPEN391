// testhps.v

// Generated using ACDS version 15.0 153

`timescale 1 ps / 1 ps
module testhps (
		input  wire        clk_clk,                         //     clk.clk
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //  hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //        .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //        .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //        .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //        .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //        .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //        .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //        .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //        .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //        .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //        .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //        .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //        .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //        .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //        .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //        .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //        .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //        .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //        .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //        .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //        .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //        .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //        .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //        .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //        .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //        .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //        .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //        .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //        .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //        .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //        .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //        .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //        .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //        .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //        .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //        .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //        .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //        .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,     //        .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //        .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //        .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //        .hps_io_i2c0_inst_SCL
		output wire [14:0] hps_mem_mem_a,                   // hps_mem.mem_a
		output wire [2:0]  hps_mem_mem_ba,                  //        .mem_ba
		output wire        hps_mem_mem_ck,                  //        .mem_ck
		output wire        hps_mem_mem_ck_n,                //        .mem_ck_n
		output wire        hps_mem_mem_cke,                 //        .mem_cke
		output wire        hps_mem_mem_cs_n,                //        .mem_cs_n
		output wire        hps_mem_mem_ras_n,               //        .mem_ras_n
		output wire        hps_mem_mem_cas_n,               //        .mem_cas_n
		output wire        hps_mem_mem_we_n,                //        .mem_we_n
		output wire        hps_mem_mem_reset_n,             //        .mem_reset_n
		inout  wire [31:0] hps_mem_mem_dq,                  //        .mem_dq
		inout  wire [3:0]  hps_mem_mem_dqs,                 //        .mem_dqs
		inout  wire [3:0]  hps_mem_mem_dqs_n,               //        .mem_dqs_n
		output wire        hps_mem_mem_odt,                 //        .mem_odt
		output wire [3:0]  hps_mem_mem_dm,                  //        .mem_dm
		input  wire        hps_mem_oct_rzqin,               //        .oct_rzqin
		input  wire        reset_reset_n,                   //   reset.reset_n
		output wire        vga_CLK,                         //     vga.CLK
		output wire        vga_HS,                          //        .HS
		output wire        vga_VS,                          //        .VS
		output wire        vga_BLANK,                       //        .BLANK
		output wire        vga_SYNC,                        //        .SYNC
		output wire [7:0]  vga_R,                           //        .R
		output wire [7:0]  vga_G,                           //        .G
		output wire [7:0]  vga_B                            //        .B
	);

	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                      // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                       // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                      // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;              // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         video_dma_controller_0_avalon_pixel_source_valid;                             // video_dma_controller_0:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [23:0] video_dma_controller_0_avalon_pixel_source_data;                              // video_dma_controller_0:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         video_dma_controller_0_avalon_pixel_source_ready;                             // video_rgb_resampler_0:stream_in_ready -> video_dma_controller_0:stream_ready
	wire         video_dma_controller_0_avalon_pixel_source_startofpacket;                     // video_dma_controller_0:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_dma_controller_0_avalon_pixel_source_endofpacket;                       // video_dma_controller_0:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                                // video_rgb_resampler_0:stream_out_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                 // video_rgb_resampler_0:stream_out_data -> video_dual_clock_buffer_0:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                                // video_dual_clock_buffer_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                        // video_rgb_resampler_0:stream_out_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                          // video_rgb_resampler_0:stream_out_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         video_pll_0_vga_clk_clk;                                                      // video_pll_0:vga_clk_clk -> [rst_controller_001:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	wire         video_dma_controller_0_avalon_dma_master_waitrequest;                         // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_waitrequest -> video_dma_controller_0:master_waitrequest
	wire  [31:0] video_dma_controller_0_avalon_dma_master_readdata;                            // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdata -> video_dma_controller_0:master_readdata
	wire  [31:0] video_dma_controller_0_avalon_dma_master_address;                             // video_dma_controller_0:master_address -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_address
	wire         video_dma_controller_0_avalon_dma_master_read;                                // video_dma_controller_0:master_read -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_read
	wire         video_dma_controller_0_avalon_dma_master_readdatavalid;                       // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_readdatavalid -> video_dma_controller_0:master_readdatavalid
	wire         video_dma_controller_0_avalon_dma_master_lock;                                // video_dma_controller_0:master_arbiterlock -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_lock
	wire   [1:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awburst;                              // mm_interconnect_0:hps_0_f2h_sdram0_data_awburst -> hps_0:f2h_sdram0_AWBURST
	wire   [3:0] mm_interconnect_0_hps_0_f2h_sdram0_data_arlen;                                // mm_interconnect_0:hps_0_f2h_sdram0_data_arlen -> hps_0:f2h_sdram0_ARLEN
	wire   [7:0] mm_interconnect_0_hps_0_f2h_sdram0_data_wstrb;                                // mm_interconnect_0:hps_0_f2h_sdram0_data_wstrb -> hps_0:f2h_sdram0_WSTRB
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_wready;                               // hps_0:f2h_sdram0_WREADY -> mm_interconnect_0:hps_0_f2h_sdram0_data_wready
	wire   [7:0] mm_interconnect_0_hps_0_f2h_sdram0_data_rid;                                  // hps_0:f2h_sdram0_RID -> mm_interconnect_0:hps_0_f2h_sdram0_data_rid
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_rready;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_rready -> hps_0:f2h_sdram0_RREADY
	wire   [3:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awlen;                                // mm_interconnect_0:hps_0_f2h_sdram0_data_awlen -> hps_0:f2h_sdram0_AWLEN
	wire   [7:0] mm_interconnect_0_hps_0_f2h_sdram0_data_wid;                                  // mm_interconnect_0:hps_0_f2h_sdram0_data_wid -> hps_0:f2h_sdram0_WID
	wire   [3:0] mm_interconnect_0_hps_0_f2h_sdram0_data_arcache;                              // mm_interconnect_0:hps_0_f2h_sdram0_data_arcache -> hps_0:f2h_sdram0_ARCACHE
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_wvalid;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_wvalid -> hps_0:f2h_sdram0_WVALID
	wire  [31:0] mm_interconnect_0_hps_0_f2h_sdram0_data_araddr;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_araddr -> hps_0:f2h_sdram0_ARADDR
	wire   [2:0] mm_interconnect_0_hps_0_f2h_sdram0_data_arprot;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_arprot -> hps_0:f2h_sdram0_ARPROT
	wire   [2:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awprot;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_awprot -> hps_0:f2h_sdram0_AWPROT
	wire  [63:0] mm_interconnect_0_hps_0_f2h_sdram0_data_wdata;                                // mm_interconnect_0:hps_0_f2h_sdram0_data_wdata -> hps_0:f2h_sdram0_WDATA
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_arvalid;                              // mm_interconnect_0:hps_0_f2h_sdram0_data_arvalid -> hps_0:f2h_sdram0_ARVALID
	wire   [3:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awcache;                              // mm_interconnect_0:hps_0_f2h_sdram0_data_awcache -> hps_0:f2h_sdram0_AWCACHE
	wire   [7:0] mm_interconnect_0_hps_0_f2h_sdram0_data_arid;                                 // mm_interconnect_0:hps_0_f2h_sdram0_data_arid -> hps_0:f2h_sdram0_ARID
	wire   [1:0] mm_interconnect_0_hps_0_f2h_sdram0_data_arlock;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_arlock -> hps_0:f2h_sdram0_ARLOCK
	wire   [1:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awlock;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_awlock -> hps_0:f2h_sdram0_AWLOCK
	wire  [31:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awaddr;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_awaddr -> hps_0:f2h_sdram0_AWADDR
	wire   [1:0] mm_interconnect_0_hps_0_f2h_sdram0_data_bresp;                                // hps_0:f2h_sdram0_BRESP -> mm_interconnect_0:hps_0_f2h_sdram0_data_bresp
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_arready;                              // hps_0:f2h_sdram0_ARREADY -> mm_interconnect_0:hps_0_f2h_sdram0_data_arready
	wire  [63:0] mm_interconnect_0_hps_0_f2h_sdram0_data_rdata;                                // hps_0:f2h_sdram0_RDATA -> mm_interconnect_0:hps_0_f2h_sdram0_data_rdata
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_awready;                              // hps_0:f2h_sdram0_AWREADY -> mm_interconnect_0:hps_0_f2h_sdram0_data_awready
	wire   [1:0] mm_interconnect_0_hps_0_f2h_sdram0_data_arburst;                              // mm_interconnect_0:hps_0_f2h_sdram0_data_arburst -> hps_0:f2h_sdram0_ARBURST
	wire   [2:0] mm_interconnect_0_hps_0_f2h_sdram0_data_arsize;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_arsize -> hps_0:f2h_sdram0_ARSIZE
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_bready;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_bready -> hps_0:f2h_sdram0_BREADY
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_rlast;                                // hps_0:f2h_sdram0_RLAST -> mm_interconnect_0:hps_0_f2h_sdram0_data_rlast
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_wlast;                                // mm_interconnect_0:hps_0_f2h_sdram0_data_wlast -> hps_0:f2h_sdram0_WLAST
	wire   [1:0] mm_interconnect_0_hps_0_f2h_sdram0_data_rresp;                                // hps_0:f2h_sdram0_RRESP -> mm_interconnect_0:hps_0_f2h_sdram0_data_rresp
	wire   [7:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awid;                                 // mm_interconnect_0:hps_0_f2h_sdram0_data_awid -> hps_0:f2h_sdram0_AWID
	wire   [7:0] mm_interconnect_0_hps_0_f2h_sdram0_data_bid;                                  // hps_0:f2h_sdram0_BID -> mm_interconnect_0:hps_0_f2h_sdram0_data_bid
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_bvalid;                               // hps_0:f2h_sdram0_BVALID -> mm_interconnect_0:hps_0_f2h_sdram0_data_bvalid
	wire   [2:0] mm_interconnect_0_hps_0_f2h_sdram0_data_awsize;                               // mm_interconnect_0:hps_0_f2h_sdram0_data_awsize -> hps_0:f2h_sdram0_AWSIZE
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_awvalid;                              // mm_interconnect_0:hps_0_f2h_sdram0_data_awvalid -> hps_0:f2h_sdram0_AWVALID
	wire         mm_interconnect_0_hps_0_f2h_sdram0_data_rvalid;                               // hps_0:f2h_sdram0_RVALID -> mm_interconnect_0:hps_0_f2h_sdram0_data_rvalid
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                              // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                                // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                                // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                               // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                                // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                                  // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                              // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                               // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                               // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                               // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                               // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                                // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                                              // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                              // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                                 // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                               // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                               // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                               // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                                              // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                                              // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                              // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                               // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                               // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                                // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                                // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                                 // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                                  // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                               // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                                              // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                               // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_readdata;   // video_dma_controller_0:slave_readdata -> mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_address;    // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_address -> video_dma_controller_0:slave_address
	wire         mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_read;       // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_read -> video_dma_controller_0:slave_read
	wire   [3:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_byteenable; // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_byteenable -> video_dma_controller_0:slave_byteenable
	wire         mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_write;      // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_write -> video_dma_controller_0:slave_write
	wire  [31:0] mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_writedata;  // mm_interconnect_1:video_dma_controller_0_avalon_dma_control_slave_writedata -> video_dma_controller_0:slave_writedata
	wire  [31:0] hps_0_f2h_irq0_irq;                                                           // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                                           // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                                               // rst_controller:reset_out -> [mm_interconnect_0:video_dma_controller_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:video_dma_controller_0_reset_reset_bridge_in_reset_reset, video_dma_controller_0:reset, video_dual_clock_buffer_0:reset_stream_in, video_rgb_resampler_0:reset]
	wire         rst_controller_001_reset_out_reset;                                           // rst_controller_001:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]
	wire         video_pll_0_reset_source_reset;                                               // video_pll_0:reset_source_reset -> rst_controller_001:reset_in0
	wire         rst_controller_002_reset_out_reset;                                           // rst_controller_002:reset_out -> [mm_interconnect_0:hps_0_f2h_sdram0_data_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire         hps_0_h2f_reset_reset;                                                        // hps_0:h2f_rst_n -> rst_controller_002:reset_in0

	testhps_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.mem_a                    (hps_mem_mem_a),                                   //            memory.mem_a
		.mem_ba                   (hps_mem_mem_ba),                                  //                  .mem_ba
		.mem_ck                   (hps_mem_mem_ck),                                  //                  .mem_ck
		.mem_ck_n                 (hps_mem_mem_ck_n),                                //                  .mem_ck_n
		.mem_cke                  (hps_mem_mem_cke),                                 //                  .mem_cke
		.mem_cs_n                 (hps_mem_mem_cs_n),                                //                  .mem_cs_n
		.mem_ras_n                (hps_mem_mem_ras_n),                               //                  .mem_ras_n
		.mem_cas_n                (hps_mem_mem_cas_n),                               //                  .mem_cas_n
		.mem_we_n                 (hps_mem_mem_we_n),                                //                  .mem_we_n
		.mem_reset_n              (hps_mem_mem_reset_n),                             //                  .mem_reset_n
		.mem_dq                   (hps_mem_mem_dq),                                  //                  .mem_dq
		.mem_dqs                  (hps_mem_mem_dqs),                                 //                  .mem_dqs
		.mem_dqs_n                (hps_mem_mem_dqs_n),                               //                  .mem_dqs_n
		.mem_odt                  (hps_mem_mem_odt),                                 //                  .mem_odt
		.mem_dm                   (hps_mem_mem_dm),                                  //                  .mem_dm
		.oct_rzqin                (hps_mem_oct_rzqin),                               //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                 //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                 //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                 //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                 //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                     //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                     //                  .hps_io_i2c0_inst_SCL
		.h2f_rst_n                (hps_0_h2f_reset_reset),                           //         h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                                         //  f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR        (mm_interconnect_0_hps_0_f2h_sdram0_data_araddr),  //   f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN         (mm_interconnect_0_hps_0_f2h_sdram0_data_arlen),   //                  .arlen
		.f2h_sdram0_ARID          (mm_interconnect_0_hps_0_f2h_sdram0_data_arid),    //                  .arid
		.f2h_sdram0_ARSIZE        (mm_interconnect_0_hps_0_f2h_sdram0_data_arsize),  //                  .arsize
		.f2h_sdram0_ARBURST       (mm_interconnect_0_hps_0_f2h_sdram0_data_arburst), //                  .arburst
		.f2h_sdram0_ARLOCK        (mm_interconnect_0_hps_0_f2h_sdram0_data_arlock),  //                  .arlock
		.f2h_sdram0_ARPROT        (mm_interconnect_0_hps_0_f2h_sdram0_data_arprot),  //                  .arprot
		.f2h_sdram0_ARVALID       (mm_interconnect_0_hps_0_f2h_sdram0_data_arvalid), //                  .arvalid
		.f2h_sdram0_ARCACHE       (mm_interconnect_0_hps_0_f2h_sdram0_data_arcache), //                  .arcache
		.f2h_sdram0_AWADDR        (mm_interconnect_0_hps_0_f2h_sdram0_data_awaddr),  //                  .awaddr
		.f2h_sdram0_AWLEN         (mm_interconnect_0_hps_0_f2h_sdram0_data_awlen),   //                  .awlen
		.f2h_sdram0_AWID          (mm_interconnect_0_hps_0_f2h_sdram0_data_awid),    //                  .awid
		.f2h_sdram0_AWSIZE        (mm_interconnect_0_hps_0_f2h_sdram0_data_awsize),  //                  .awsize
		.f2h_sdram0_AWBURST       (mm_interconnect_0_hps_0_f2h_sdram0_data_awburst), //                  .awburst
		.f2h_sdram0_AWLOCK        (mm_interconnect_0_hps_0_f2h_sdram0_data_awlock),  //                  .awlock
		.f2h_sdram0_AWPROT        (mm_interconnect_0_hps_0_f2h_sdram0_data_awprot),  //                  .awprot
		.f2h_sdram0_AWVALID       (mm_interconnect_0_hps_0_f2h_sdram0_data_awvalid), //                  .awvalid
		.f2h_sdram0_AWCACHE       (mm_interconnect_0_hps_0_f2h_sdram0_data_awcache), //                  .awcache
		.f2h_sdram0_BRESP         (mm_interconnect_0_hps_0_f2h_sdram0_data_bresp),   //                  .bresp
		.f2h_sdram0_BID           (mm_interconnect_0_hps_0_f2h_sdram0_data_bid),     //                  .bid
		.f2h_sdram0_BVALID        (mm_interconnect_0_hps_0_f2h_sdram0_data_bvalid),  //                  .bvalid
		.f2h_sdram0_BREADY        (mm_interconnect_0_hps_0_f2h_sdram0_data_bready),  //                  .bready
		.f2h_sdram0_ARREADY       (mm_interconnect_0_hps_0_f2h_sdram0_data_arready), //                  .arready
		.f2h_sdram0_AWREADY       (mm_interconnect_0_hps_0_f2h_sdram0_data_awready), //                  .awready
		.f2h_sdram0_RREADY        (mm_interconnect_0_hps_0_f2h_sdram0_data_rready),  //                  .rready
		.f2h_sdram0_RDATA         (mm_interconnect_0_hps_0_f2h_sdram0_data_rdata),   //                  .rdata
		.f2h_sdram0_RRESP         (mm_interconnect_0_hps_0_f2h_sdram0_data_rresp),   //                  .rresp
		.f2h_sdram0_RLAST         (mm_interconnect_0_hps_0_f2h_sdram0_data_rlast),   //                  .rlast
		.f2h_sdram0_RID           (mm_interconnect_0_hps_0_f2h_sdram0_data_rid),     //                  .rid
		.f2h_sdram0_RVALID        (mm_interconnect_0_hps_0_f2h_sdram0_data_rvalid),  //                  .rvalid
		.f2h_sdram0_WLAST         (mm_interconnect_0_hps_0_f2h_sdram0_data_wlast),   //                  .wlast
		.f2h_sdram0_WVALID        (mm_interconnect_0_hps_0_f2h_sdram0_data_wvalid),  //                  .wvalid
		.f2h_sdram0_WDATA         (mm_interconnect_0_hps_0_f2h_sdram0_data_wdata),   //                  .wdata
		.f2h_sdram0_WSTRB         (mm_interconnect_0_hps_0_f2h_sdram0_data_wstrb),   //                  .wstrb
		.f2h_sdram0_WREADY        (mm_interconnect_0_hps_0_f2h_sdram0_data_wready),  //                  .wready
		.f2h_sdram0_WID           (mm_interconnect_0_hps_0_f2h_sdram0_data_wid),     //                  .wid
		.h2f_axi_clk              (clk_clk),                                         //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                                //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                                //                  .awaddr
		.h2f_AWLEN                (),                                                //                  .awlen
		.h2f_AWSIZE               (),                                                //                  .awsize
		.h2f_AWBURST              (),                                                //                  .awburst
		.h2f_AWLOCK               (),                                                //                  .awlock
		.h2f_AWCACHE              (),                                                //                  .awcache
		.h2f_AWPROT               (),                                                //                  .awprot
		.h2f_AWVALID              (),                                                //                  .awvalid
		.h2f_AWREADY              (),                                                //                  .awready
		.h2f_WID                  (),                                                //                  .wid
		.h2f_WDATA                (),                                                //                  .wdata
		.h2f_WSTRB                (),                                                //                  .wstrb
		.h2f_WLAST                (),                                                //                  .wlast
		.h2f_WVALID               (),                                                //                  .wvalid
		.h2f_WREADY               (),                                                //                  .wready
		.h2f_BID                  (),                                                //                  .bid
		.h2f_BRESP                (),                                                //                  .bresp
		.h2f_BVALID               (),                                                //                  .bvalid
		.h2f_BREADY               (),                                                //                  .bready
		.h2f_ARID                 (),                                                //                  .arid
		.h2f_ARADDR               (),                                                //                  .araddr
		.h2f_ARLEN                (),                                                //                  .arlen
		.h2f_ARSIZE               (),                                                //                  .arsize
		.h2f_ARBURST              (),                                                //                  .arburst
		.h2f_ARLOCK               (),                                                //                  .arlock
		.h2f_ARCACHE              (),                                                //                  .arcache
		.h2f_ARPROT               (),                                                //                  .arprot
		.h2f_ARVALID              (),                                                //                  .arvalid
		.h2f_ARREADY              (),                                                //                  .arready
		.h2f_RID                  (),                                                //                  .rid
		.h2f_RDATA                (),                                                //                  .rdata
		.h2f_RRESP                (),                                                //                  .rresp
		.h2f_RLAST                (),                                                //                  .rlast
		.h2f_RVALID               (),                                                //                  .rvalid
		.h2f_RREADY               (),                                                //                  .rready
		.f2h_axi_clk              (clk_clk),                                         //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                                //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                                //                  .awaddr
		.f2h_AWLEN                (),                                                //                  .awlen
		.f2h_AWSIZE               (),                                                //                  .awsize
		.f2h_AWBURST              (),                                                //                  .awburst
		.f2h_AWLOCK               (),                                                //                  .awlock
		.f2h_AWCACHE              (),                                                //                  .awcache
		.f2h_AWPROT               (),                                                //                  .awprot
		.f2h_AWVALID              (),                                                //                  .awvalid
		.f2h_AWREADY              (),                                                //                  .awready
		.f2h_AWUSER               (),                                                //                  .awuser
		.f2h_WID                  (),                                                //                  .wid
		.f2h_WDATA                (),                                                //                  .wdata
		.f2h_WSTRB                (),                                                //                  .wstrb
		.f2h_WLAST                (),                                                //                  .wlast
		.f2h_WVALID               (),                                                //                  .wvalid
		.f2h_WREADY               (),                                                //                  .wready
		.f2h_BID                  (),                                                //                  .bid
		.f2h_BRESP                (),                                                //                  .bresp
		.f2h_BVALID               (),                                                //                  .bvalid
		.f2h_BREADY               (),                                                //                  .bready
		.f2h_ARID                 (),                                                //                  .arid
		.f2h_ARADDR               (),                                                //                  .araddr
		.f2h_ARLEN                (),                                                //                  .arlen
		.f2h_ARSIZE               (),                                                //                  .arsize
		.f2h_ARBURST              (),                                                //                  .arburst
		.f2h_ARLOCK               (),                                                //                  .arlock
		.f2h_ARCACHE              (),                                                //                  .arcache
		.f2h_ARPROT               (),                                                //                  .arprot
		.f2h_ARVALID              (),                                                //                  .arvalid
		.f2h_ARREADY              (),                                                //                  .arready
		.f2h_ARUSER               (),                                                //                  .aruser
		.f2h_RID                  (),                                                //                  .rid
		.f2h_RDATA                (),                                                //                  .rdata
		.f2h_RRESP                (),                                                //                  .rresp
		.f2h_RLAST                (),                                                //                  .rlast
		.f2h_RVALID               (),                                                //                  .rvalid
		.f2h_RREADY               (),                                                //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                 //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                 //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                 //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                 //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                 //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                 //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                 //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                 //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                  //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                              //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                               //          f2h_irq1.irq
	);

	testhps_video_dma_controller_0 video_dma_controller_0 (
		.clk                  (clk_clk),                                                                      //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                                               //                    reset.reset
		.master_address       (video_dma_controller_0_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma_controller_0_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_arbiterlock   (video_dma_controller_0_avalon_dma_master_lock),                                //                         .lock
		.master_read          (video_dma_controller_0_avalon_dma_master_read),                                //                         .read
		.master_readdata      (video_dma_controller_0_avalon_dma_master_readdata),                            //                         .readdata
		.master_readdatavalid (video_dma_controller_0_avalon_dma_master_readdatavalid),                       //                         .readdatavalid
		.slave_address        (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                         .readdata
		.stream_ready         (video_dma_controller_0_avalon_pixel_source_ready),                             //      avalon_pixel_source.ready
		.stream_data          (video_dma_controller_0_avalon_pixel_source_data),                              //                         .data
		.stream_startofpacket (video_dma_controller_0_avalon_pixel_source_startofpacket),                     //                         .startofpacket
		.stream_endofpacket   (video_dma_controller_0_avalon_pixel_source_endofpacket),                       //                         .endofpacket
		.stream_valid         (video_dma_controller_0_avalon_pixel_source_valid)                              //                         .valid
	);

	testhps_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (clk_clk),                                                         //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                                  //         reset_stream_in.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                                         //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_001_reset_out_reset),                              //        reset_stream_out.reset
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),                   //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket),           //                        .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),             //                        .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),                   //                        .valid
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),                    //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	testhps_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),                 //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)  // reset_source.reset
	);

	testhps_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clk_clk),                                                  //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                           //             reset.reset
		.stream_in_startofpacket  (video_dma_controller_0_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_dma_controller_0_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_dma_controller_0_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (video_dma_controller_0_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (video_dma_controller_0_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),            // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),    //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),      //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),            //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)              //                  .data
	);

	testhps_video_vga_controller_0 video_vga_controller_0 (
		.clk           (video_pll_0_vga_clk_clk),                                         //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),                              //              reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_CLK),                                                         // external_interface.export
		.VGA_HS        (vga_HS),                                                          //                   .export
		.VGA_VS        (vga_VS),                                                          //                   .export
		.VGA_BLANK     (vga_BLANK),                                                       //                   .export
		.VGA_SYNC      (vga_SYNC),                                                        //                   .export
		.VGA_R         (vga_R),                                                           //                   .export
		.VGA_G         (vga_G),                                                           //                   .export
		.VGA_B         (vga_B)                                                            //                   .export
	);

	testhps_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_sdram0_data_awid                                         (mm_interconnect_0_hps_0_f2h_sdram0_data_awid),           //                                        hps_0_f2h_sdram0_data.awid
		.hps_0_f2h_sdram0_data_awaddr                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_awaddr),         //                                                             .awaddr
		.hps_0_f2h_sdram0_data_awlen                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_awlen),          //                                                             .awlen
		.hps_0_f2h_sdram0_data_awsize                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_awsize),         //                                                             .awsize
		.hps_0_f2h_sdram0_data_awburst                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_awburst),        //                                                             .awburst
		.hps_0_f2h_sdram0_data_awlock                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_awlock),         //                                                             .awlock
		.hps_0_f2h_sdram0_data_awcache                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_awcache),        //                                                             .awcache
		.hps_0_f2h_sdram0_data_awprot                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_awprot),         //                                                             .awprot
		.hps_0_f2h_sdram0_data_awvalid                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_awvalid),        //                                                             .awvalid
		.hps_0_f2h_sdram0_data_awready                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_awready),        //                                                             .awready
		.hps_0_f2h_sdram0_data_wid                                          (mm_interconnect_0_hps_0_f2h_sdram0_data_wid),            //                                                             .wid
		.hps_0_f2h_sdram0_data_wdata                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_wdata),          //                                                             .wdata
		.hps_0_f2h_sdram0_data_wstrb                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_wstrb),          //                                                             .wstrb
		.hps_0_f2h_sdram0_data_wlast                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_wlast),          //                                                             .wlast
		.hps_0_f2h_sdram0_data_wvalid                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_wvalid),         //                                                             .wvalid
		.hps_0_f2h_sdram0_data_wready                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_wready),         //                                                             .wready
		.hps_0_f2h_sdram0_data_bid                                          (mm_interconnect_0_hps_0_f2h_sdram0_data_bid),            //                                                             .bid
		.hps_0_f2h_sdram0_data_bresp                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_bresp),          //                                                             .bresp
		.hps_0_f2h_sdram0_data_bvalid                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_bvalid),         //                                                             .bvalid
		.hps_0_f2h_sdram0_data_bready                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_bready),         //                                                             .bready
		.hps_0_f2h_sdram0_data_arid                                         (mm_interconnect_0_hps_0_f2h_sdram0_data_arid),           //                                                             .arid
		.hps_0_f2h_sdram0_data_araddr                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_araddr),         //                                                             .araddr
		.hps_0_f2h_sdram0_data_arlen                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_arlen),          //                                                             .arlen
		.hps_0_f2h_sdram0_data_arsize                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_arsize),         //                                                             .arsize
		.hps_0_f2h_sdram0_data_arburst                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_arburst),        //                                                             .arburst
		.hps_0_f2h_sdram0_data_arlock                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_arlock),         //                                                             .arlock
		.hps_0_f2h_sdram0_data_arcache                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_arcache),        //                                                             .arcache
		.hps_0_f2h_sdram0_data_arprot                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_arprot),         //                                                             .arprot
		.hps_0_f2h_sdram0_data_arvalid                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_arvalid),        //                                                             .arvalid
		.hps_0_f2h_sdram0_data_arready                                      (mm_interconnect_0_hps_0_f2h_sdram0_data_arready),        //                                                             .arready
		.hps_0_f2h_sdram0_data_rid                                          (mm_interconnect_0_hps_0_f2h_sdram0_data_rid),            //                                                             .rid
		.hps_0_f2h_sdram0_data_rdata                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_rdata),          //                                                             .rdata
		.hps_0_f2h_sdram0_data_rresp                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_rresp),          //                                                             .rresp
		.hps_0_f2h_sdram0_data_rlast                                        (mm_interconnect_0_hps_0_f2h_sdram0_data_rlast),          //                                                             .rlast
		.hps_0_f2h_sdram0_data_rvalid                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_rvalid),         //                                                             .rvalid
		.hps_0_f2h_sdram0_data_rready                                       (mm_interconnect_0_hps_0_f2h_sdram0_data_rready),         //                                                             .rready
		.clk_0_clk_clk                                                      (clk_clk),                                                //                                                    clk_0_clk.clk
		.hps_0_f2h_sdram0_data_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                     // hps_0_f2h_sdram0_data_agent_reset_sink_reset_bridge_in_reset.reset
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                         //           video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_avalon_dma_master_address                   (video_dma_controller_0_avalon_dma_master_address),       //                     video_dma_controller_0_avalon_dma_master.address
		.video_dma_controller_0_avalon_dma_master_waitrequest               (video_dma_controller_0_avalon_dma_master_waitrequest),   //                                                             .waitrequest
		.video_dma_controller_0_avalon_dma_master_read                      (video_dma_controller_0_avalon_dma_master_read),          //                                                             .read
		.video_dma_controller_0_avalon_dma_master_readdata                  (video_dma_controller_0_avalon_dma_master_readdata),      //                                                             .readdata
		.video_dma_controller_0_avalon_dma_master_readdatavalid             (video_dma_controller_0_avalon_dma_master_readdatavalid), //                                                             .readdatavalid
		.video_dma_controller_0_avalon_dma_master_lock                      (video_dma_controller_0_avalon_dma_master_lock)           //                                                             .lock
	);

	testhps_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                                 //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                               //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                                //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                               //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                                              //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                               //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                                              //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                               //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                                              //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                                              //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                                  //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                                //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                                //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                                //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                               //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                               //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                                  //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                                //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                               //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                               //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                                 //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                               //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                                //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                               //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                                              //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                               //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                                              //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                               //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                                              //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                                              //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                                  //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                                //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                                //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                                //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                               //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                               //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                                      //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                           // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                               //            video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_avalon_dma_control_slave_address             (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_address),    //               video_dma_controller_0_avalon_dma_control_slave.address
		.video_dma_controller_0_avalon_dma_control_slave_write               (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_write),      //                                                              .write
		.video_dma_controller_0_avalon_dma_control_slave_read                (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_read),       //                                                              .read
		.video_dma_controller_0_avalon_dma_control_slave_readdata            (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                                                              .readdata
		.video_dma_controller_0_avalon_dma_control_slave_writedata           (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                                                              .writedata
		.video_dma_controller_0_avalon_dma_control_slave_byteenable          (mm_interconnect_1_video_dma_controller_0_avalon_dma_control_slave_byteenable)  //                                                              .byteenable
	);

	testhps_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	testhps_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
